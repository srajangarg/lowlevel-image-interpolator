--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   01:03:31 04/06/2016
-- Design Name:   
-- Module Name:   /home/anuj/DLDProject/ImageInterpolator/test2.vhd
-- Project Name:  ImageInterpolator
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: interpolator_top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY test2 IS
END test2;
 
ARCHITECTURE behavior OF test2 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT interpolator_top
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         start : IN  std_logic;
         RPixel : IN  std_logic_vector(15 downto 0);
         GPixel : IN  std_logic_vector(15 downto 0);
         BPixel : IN  std_logic_vector(15 downto 0);
         outRPixel : INOUT  std_logic_vector(15 downto 0);
         outGPixel : INOUT  std_logic_vector(15 downto 0);
         outBPixel : INOUT  std_logic_vector(15 downto 0);
         outputReady : INOUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal start : std_logic := '0';
   signal RPixel : std_logic_vector(15 downto 0) := (others => '0');
   signal GPixel : std_logic_vector(15 downto 0) := (others => '0');
   signal BPixel : std_logic_vector(15 downto 0) := (others => '0');

	--BiDirs
   signal outRPixel : std_logic_vector(15 downto 0);
   signal outGPixel : std_logic_vector(15 downto 0);
   signal outBPixel : std_logic_vector(15 downto 0);
   signal outputReady : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: interpolator_top PORT MAP (
          clk => clk,
          reset => reset,
          start => start,
          RPixel => RPixel,
          GPixel => GPixel,
          BPixel => BPixel,
          outRPixel => outRPixel,
          outGPixel => outGPixel,
          outBPixel => outBPixel,
          outputReady => outputReady
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
    reset<='1';
    wait for clk_period*5;
    reset<='0';
     start<='1';
    RPixel <= "1000000000000000";
    GPixel <= "1000000000000000";
    BPixel <= "1000000000000000";
    wait for clk_period*2;
    start<='0';
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011100101";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111001";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111100";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111100";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011101110";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011110101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111110";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011111010";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000011001100";
    BPixel<="0000000010111101";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001100000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000101111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000101000";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001000100";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001110110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011011001";
    BPixel<="0000000011000111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011110001";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011110110";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111011";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110110";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011110010";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011110000";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011110010";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111011";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011110010";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110101";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110111";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011111000";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111110";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111001";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011101101";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011101000";
    BPixel<="0000000011010101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101110";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011100011";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011101110";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101111";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111010";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110001";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010101110";
    BPixel<="0000000010101001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000111000";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000001000101";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001101001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010010110";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110111";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010011001";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001010000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000000101010";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010111010";
    BPixel<="0000000010011011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011111011";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011101110";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110111";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110011";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110101";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110010";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110001";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011101011";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010011100";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001010010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001011000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000110101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001010110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000010100010";
    BPixel<="0000000010011000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000011000011";
    BPixel<="0000000010011111";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000010001101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011011001";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001101";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101011";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000110";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011100101";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011001000";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001100001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010110011";
    BPixel<="0000000010110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011100001";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011101110";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011110101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011101001";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000010000111";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000110101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000001000001";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000001011110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000010100011";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111110";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111000";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110011";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111000";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111010";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101110";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110001";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001001011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001011010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001111011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001100111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001000110";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000011011";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010101110";
    BPixel<="0000000010011001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100100";
    BPixel<="0000000011011001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010010000";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001001111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001100111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010110101";
    BPixel<="0000000010100010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011100110";
    BPixel<="0000000011011001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000101000";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001011110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011011101";
    BPixel<="0000000010001010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011001011";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010111001";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011011010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000010001110";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000010000000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000001001000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101110";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101010";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000010001111";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000001000111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000010000110";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001100010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001000111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011011100";
    BPixel<="0000000011001101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110101";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011100101";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101010";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011101011";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001011110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000001001100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011011100";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000010011011";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001100";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011110";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011000";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010010101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010000010";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010111011";
    BPixel<="0000000010101000";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011011010";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011010001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011010001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000110";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010111001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001111";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010011111";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010110001";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000111011";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000100010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001100";
    BPixel<="0000000011000000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001000";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001111101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011001111";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011000001";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010100110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001010";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101011";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001001100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011101110";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101001";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011110001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111101";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110010";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110010";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110011";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010010011";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010110011";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111100";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010101100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101101";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001011101";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001000100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001001010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001011110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010101000";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000101";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010010";
    BPixel<="0000000001111101";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010100000";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001000001";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001111011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010111";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011001001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011100001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101001";
    BPixel<="0000000001111100";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001100111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011010111";
    BPixel<="0000000011000100";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000101101";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010001011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000111";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010110100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011001000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011100010";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010110110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000100010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011011100";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111101";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111100";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011101101";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101001";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010011000";
    BPixel<="0000000010100000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000111010";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000010010111";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000011000100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000110";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011011010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010101101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010000";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000001000100";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001111010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001011000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010001010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011100000";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000011000110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011011001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011010101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000101";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010111000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010111000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001001000";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000010";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010101001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010111101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010110100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101110";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010111101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010110010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000010110100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010011010";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001010";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001111110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000100011";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011101000";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111011";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110011";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111010";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011000110";
    BPixel<="0000000010110000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000010001110";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001101011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001111011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000010100100";
    BPixel<="0000000010000000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011011010";
    BPixel<="0000000010111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011100110";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010111010";
    BPixel<="0000000010101011";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010111010";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111010";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011000101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010100100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010101111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011011001";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000001001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001000";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010101000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010101000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011000010";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010001100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111110";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010010";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011000101";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011101010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011010000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011111";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000010010010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000111010";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010100101";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010110110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001100";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011100";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011011110";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011010010";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010001010";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111000";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011101100";
    BPixel<="0000000011011110";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010001110";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000001010100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001100111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001111001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010111010";
    BPixel<="0000000010011011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011100100";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000010010010";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000101111";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101100";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011010000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011010101";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010001";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001101";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001111";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010100100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001101101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000010000010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011011101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011000111";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011101000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011001101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011001101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010001";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001010111";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000101";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111110";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111001";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010000000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011000010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010110111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000010110011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010110010";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110001";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111010";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001000101";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010001010";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110010";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010000";
    BPixel<="0000000011000001";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000001001110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000110011";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001011101";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001011101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000111100";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000101001";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010100101";
    BPixel<="0000000010001011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011100110";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011110000";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011110000";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011001001";
    BPixel<="0000000010110001";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000010000000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111011";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111110";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010110101";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110011";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000001001010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000001101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000101";
    BPixel<="0000000010101101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010011111";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111110";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010111110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000010110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010011111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011110";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010010100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010101001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111010";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110111";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001010011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001010010";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011001110";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011001100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010110";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011001011";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011010011";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011010110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011100001";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001011111";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010010110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000000";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011011000";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010100";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011011111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011000110";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000001000001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001010";
    BPixel<="0000000010111100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000010010110";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000001000011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001100000";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001110101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000010001111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000110011";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010111101";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110011";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110010";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110011";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011010101";
    BPixel<="0000000011000101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000100101";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000010010000";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110011";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011011000";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011100011";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011101001";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000011001010";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000010001011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000101010";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001000101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000010010011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011100010";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010001";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011001111";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001110";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010111100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010110000";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000001001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010011";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000111";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010101111";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010100111";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010011101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010010101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010010110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010010101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010011000";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001001110";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001001011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010001000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010010101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010101111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010100110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010011000";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000110010";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010100010";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011100";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001111";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010110110";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010101110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010101001";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010110100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011000101";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001000011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001101100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000010000011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000101";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010101000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010110011";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000111";
    BPixel<="0000000010001011";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001010001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001011110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110010";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110010";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111001";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011100100";
    BPixel<="0000000011010000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010100001";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110110";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010101110";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101101";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010011001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011000";
    BPixel<="0000000010001100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010001100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000000000110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011000011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010101000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010110000";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010101110";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010011101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000010001101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001100001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001000101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000000111000";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000000101011";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001000111";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001100010";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010010010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010000111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000010110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001101100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011011001";
    BPixel<="0000000010000010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011100000";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011100010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001100000";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001011111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000101";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011100010";
    BPixel<="0000000010000000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011001000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011001010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011010001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011001111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011010000";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011100001";
    BPixel<="0000000010011001";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000110010";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010100110";
    BPixel<="0000000010011001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011101100";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000001100001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001110001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110001";
    BPixel<="0000000010011101";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011010000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011100001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010010";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010100";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010011";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001111001";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000010100010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010110010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010011";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110011";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010000111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001010001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000000111011";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001110100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001110100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001111110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001111000";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001001010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001000110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000000111111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000000110011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000101100";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000000111110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010001101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111101";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010111111";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111001";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010010001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001101010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001111";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010001000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011001000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010100111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010101111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011000001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000000";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000010010001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000011001001";
    BPixel<="0000000010101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110010";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111110";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000011000110";
    BPixel<="0000000010101001";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010100100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001001";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010100100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010101010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010110100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010101100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010110111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011001000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010100000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001111101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111011";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001111111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000111110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000001";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111001";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110011";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010000001";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010000110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001111111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001011000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001001001";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001101001";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010110110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011001110";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010111101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000111100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001111011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011010";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011011010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001010";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011000100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011101001";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001111111";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110101";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111001";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010011001";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000111101";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011100100";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111111";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000010";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011001101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011010011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011011011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010110011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000001001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111011";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111111";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001000100";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010000111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001100110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001111000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001111000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100110";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001100110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001010101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000111000";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000101011";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001001011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000111010";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001100";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010100101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000001";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010100110";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011000001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000010000000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000001000001";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111000";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110001";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011011000";
    BPixel<="0000000010111110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011100111";
    BPixel<="0000000010111101";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001011100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001010010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011000";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010100011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010011110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011000110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110101";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000101";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001100111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000000110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000000111011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001100110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001101101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001111000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001000010";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001010010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010011111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001110";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011010";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110111";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011001100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011010100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010111010";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011011101";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011101011";
    BPixel<="0000000011010110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010110000";
    BPixel<="0000000010011100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000010011111";
    BPixel<="0000000010001100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000010011000";
    BPixel<="0000000010000101";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010110001";
    BPixel<="0000000010100000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011011111";
    BPixel<="0000000011010000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111110";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001111000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001010110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000000110111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000111100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010100001";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001011100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001011010";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011111";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011000111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011000000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011011111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010111000";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000001";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010000111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010010011";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001111";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001000111";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010011010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000000";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010010100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010110111";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001110101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000101101";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000100100";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000010001100";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011110001";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011101111";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110011";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111101";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111011";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001110011";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010011000";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010001111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010011110";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001111010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001100110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010011101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010000101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000010010000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010011001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001101110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001101110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010000100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010001001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010001100";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001111111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011001111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011110";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010000010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011101001";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010100000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000000000100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000111001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000001000000";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001110010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010111000";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010011";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001101";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110011";
    BPixel<="0000000010010100";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011010010";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000010101001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001000010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110111";
    BPixel<="0000000011011110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111011";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010100001";
    BPixel<="0000000010011111";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000111111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011011011";
    BPixel<="0000000010011000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011100011";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011000111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011001101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011010111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101101";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010100";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000010001011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000001000100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010100000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011100100";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011001";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010100111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010010000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010001111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010010101";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010011011";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001111001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001111101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001101111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001101110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000010010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001100000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000001";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110010";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000010001001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000111100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010011011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010100101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111100";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110001";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111001";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000010011000";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000100000";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000011010101";
    BPixel<="0000000010111111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011111010";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011111101";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011101101";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010001110";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000001000101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011001100";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111000";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010011110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011000101";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010110001";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001011010";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001100101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001110011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001100010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010010101";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010010111";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010000010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011001010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011011000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011011101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000010010110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001101111";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011100000";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011101010";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011000011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011011010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011100000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010111110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101010";
    BPixel<="0000000010011010";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001011000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001100001";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001100001";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001111110";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011101101";
    BPixel<="0000000010001011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011011000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001110";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010010";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001110110";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010101111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001010";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001001";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000000111100";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010001000";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010010110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010000000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001111101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001101111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111001";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010100101";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010110100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010111110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010100110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101111";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001010001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001110110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010011111";
    BPixel<="0000000010010011";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001011";
    BPixel<="0000000010001010";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101101";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010110011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010110101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010101110";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010111100";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001000010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000100011";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001011111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010000111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010000010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010010101";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010011110";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000001";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000110111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110011";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010011111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001110";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011001101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011011010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011100000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001000";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001100";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011100101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011001000";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011010011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101011";
    BPixel<="0000000010000000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000001001011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001111011";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000011000001";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011010111";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011100100";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000111";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010011";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011011001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011001";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000111";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001001110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001000011";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001000011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000101101";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010010011";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010001101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010001000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010001010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000001111110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001101111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001001001";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000011111";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000110110";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010110110";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010001111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011000001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001000";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001101110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000101110";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011011";
    BPixel<="0000000011010111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110011";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111000";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011101110";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010000111";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010000010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001011";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011000110";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001001110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000101011";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100100";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001000011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010000000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000001111100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000001111111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010001110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010010000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010011011";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000000011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010010100";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000110";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011100000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010101110";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011000110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011001111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011011101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011010";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010011001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000001000111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110001";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011101001";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110000";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000010000010";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011100";
    BPixel<="0000000010000000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010111101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010101110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010100000";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010000";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010100010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010000010";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010001100";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010000010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111011";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010000011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010000111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111100";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010000011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001111010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001101110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001010111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110100";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111011";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110111";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001100000";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001011101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001001011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000101101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001011101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000001010000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010101111";
    BPixel<="0000000010011001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110010";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111011";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000111111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001101011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001011110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010000101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001110100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001011010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001001110";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000000001001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000010010100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001110000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001010001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001111001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001101011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001110001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001111001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001110000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001110000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010000001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010000000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010000001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000011";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000111";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001110011";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001000011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011010011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011000011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011100010";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010001111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000001000110";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110100";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110001";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011101010";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011101100";
    BPixel<="0000000011011110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111010";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110011";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011011110";
    BPixel<="0000000010111111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010110011";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001101011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001110100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001010110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000001000011";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000100110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010011100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011100101";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011000010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011011001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011010101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011010101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101110";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010001001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010001111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010001010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001111011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000111011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000111001";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001010001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001110110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010000100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001011000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001000111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001101010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100001";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011111";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011011";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001011001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001100101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001000110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001111100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010100111";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110001";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000001";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000010";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111111";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000101";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001101";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010011011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001101110";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011110111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111001";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100100";
    BPixel<="0000000011010100";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010010100";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000111";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010100011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010010111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010101001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001010";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010111100";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010010011";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001010101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001011010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001011110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011100";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011011";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001111010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001011111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000100000";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000010110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000110010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111110";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001010000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000101000";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000000111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000110000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001101110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010000000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001111011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010001110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010001111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010001011";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001000111";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011100010";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010111";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000010000100";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001000001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001011001";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001110101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001110011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001011001";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001101101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011101101";
    BPixel<="0000000011010011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111000";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000011000000";
    BPixel<="0000000010111101";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000001001110";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010110111";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011011100";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011011110";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011100011";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011110";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010111010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000110111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100111";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000100";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010000110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010001111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010000010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010000011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010000001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010000100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110001";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000101001";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000101001";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000101001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000011000";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000100011";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001111001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010000001";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001000100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000101001";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000010011";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000000010101";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000101110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010000001";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001011110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001001101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001100010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000000111101";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001010011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111001";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111110";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010010011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010101000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110000";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101110";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000100111";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011010110";
    BPixel<="0000000011001011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110100";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100001";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000101100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001111000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111011";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010100110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101000";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010111011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001101111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001111110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001000101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001011001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001111110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000010111";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000010011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000101001";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011011111";
    BPixel<="0000000011010010";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001101000";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000111010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001110010";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011101";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000010101";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000000011000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001101111";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011011101";
    BPixel<="0000000011001111";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001110001";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001111101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111000";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010001100";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110110";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010000000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110111";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010100100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011011110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011100010";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010111111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011100000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101011";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011101110";
    BPixel<="0000000010001100";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001111001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000100101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011010000";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001101010";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000111011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000010101011";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011001010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011001001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011011100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011001";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010001111";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000111110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010001000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110010";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010001010";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010010001";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000001111110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000001111100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010001000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000111101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000010000011";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001101001";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000000001100";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000100101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000011101";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001101001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001111010";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000110011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000010001110";
    BPixel<="0000000001111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000100110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000010011";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000010101";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001111001";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001010101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001001000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001010111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010101";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010101100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010101100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000010111011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011000111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110111";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000111101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001100100";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110000";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110000";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011100";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000010111";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001011011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000001";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110011";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011110";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001001110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001000110";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001001100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001010111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001010101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001111000";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000000000110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000101011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000011011";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000101000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000101000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000110100";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001011111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010001000";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001101000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000000000111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000110000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000011101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000101001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001101010";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000111010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000100010";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010000100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010000011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000001111110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000001111100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010000011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010000111";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000000111110";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000110010";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001000010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000010010001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011000010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011010011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011011010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001110";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011101110";
    BPixel<="0000000010001000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010100100";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000100110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000100100";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010110011";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011100110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011000101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011011110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011010100";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011010010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011010100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010010";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011001011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000010";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010000000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010000010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000001111101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010000000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001001111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000110001";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000001111";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000000010011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000000011010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000000100011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000100100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000011001";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001100110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010001010";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000111101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000001110";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000010000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000011000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000010110";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011010";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001111000";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001101101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001010101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001010111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001010011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001000110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010001111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110010";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010101100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010111010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010111100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001101111";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000010101000";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101110";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011011100";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011101010";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010111001";
    BPixel<="0000000001111101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000001000000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010100011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010100";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110110";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001011100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001001111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001010101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001010111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001101101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001110111";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011101";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000011100";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000011011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010101";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000001000001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010001010";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001100000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000011111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000000100011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000000100001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000011111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000010010";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000110011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001001111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001101111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001111100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001000111";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010110001";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011001000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011001011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011001100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011010100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011101011";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000010011011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000110110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001101110";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000001000010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000010011111";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011010010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011100001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010100";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001000";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011010101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011010001";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010110";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001001";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010001111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001111100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000110110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000000010111";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000100011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000100011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000000100010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000000011101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010001010";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000001000001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010110";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000011001";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000100000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000011000";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001110100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001010110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001010011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001001100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010111";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001110";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001010000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000101011";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010010110";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001010101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000001001100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001000011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000001000010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001110000";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011001011";
    BPixel<="0000000010110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110011";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101000";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000010011000";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000100110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000111011";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001110010";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001100110";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001101001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010000010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001011000";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000100100";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001110";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001101";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010000";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001111";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001001111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001010101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001010110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001110101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000010011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000011000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000010011";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000010011";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001000000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010001010";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001100100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000010111";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000000100001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000000100010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000011100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000011010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000111001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001111010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010000101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000110101";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011100000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001010";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011001";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010111111";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000110100";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000011000110";
    BPixel<="0000000010111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001101010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000111011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101011";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011011011";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011001011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011011010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011011011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011001101";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011100011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011010010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011000110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010101001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111100";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000001111100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001111001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001111000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001001110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000110101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000010111";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000011111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000000100010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000000100010";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000010111";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001100101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010001011";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000001000010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000010111";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011000";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000010101";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001110101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001010101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001010001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001001101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001000010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001001000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000110100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000101100";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010010010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111101";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000001";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001001";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010101100";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011000111";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000010000000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010111010";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000001001101";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001110010";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011100110";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010111000";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010101000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010101000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010110000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010101110";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000110100";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001001111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001000100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001000111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001001110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001110010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000010101";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000100000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000011101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000011000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001000000";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001010110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010001010";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001100010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000000010010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000011100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000000100001";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000100101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000100111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000000010100";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000110011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001101101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001111000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001110111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000001111011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001111101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010010001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011000110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010001";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011011110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011010010";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011000100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011100010";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001010000";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000001000011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011110011";
    BPixel<="0000000011001110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110110";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011011100";
    BPixel<="0000000010111101";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000110110";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000001000100";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010100001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110001";
    BPixel<="0000000010001010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000110";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011010010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001101100";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010001000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000001111100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001110101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001101110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000110101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000010111";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000100101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000100010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000011111";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000011100";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010001011";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001000011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000011001";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000011001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000011011";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010100";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001111011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001010101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001010010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001010000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010100";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101000";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010110111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010100111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011000111";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010110100";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010100001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010111111";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011000010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101110";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101000";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011000110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010001001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000000111111";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010100";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001100";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011100";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001010011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001010101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010001";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010001111";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000100111";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000010111";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000011000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000010101";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000011011";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001001111";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010001100";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000100001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000011110";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000011010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000000011001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000011011";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000000111011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001101111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010000100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001111000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010000110";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010000101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001001100";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010110000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011010011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011100000";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010010";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001100";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001011111";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011110010";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011110111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011100110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010101011";
    BPixel<="0000000010001110";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000001000010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001101011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010100000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011000011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011000";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010100";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111001";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000111101";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010000000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001111000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001101101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000111010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000110010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000010101";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000100001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000011000";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000111000";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010000101";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001100001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000001000001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000000011100";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000010011";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000101110";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001010110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001000101";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001010101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010010101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011000010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110010";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110111";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101100";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011101000";
    BPixel<="0000000010011011";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000001000011";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001110110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010111110";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001100101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001101";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010110011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010101001";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010011110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001001101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010100";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000000111100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010111";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001100101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001010010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001100010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001001101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000101011";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000100000";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000100011";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001010101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000001110110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000001110110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000000110111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001101110";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000001000010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000111101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001000110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000001000101";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000110001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001000111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010101001";
    BPixel<="0000000010110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011101000";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001100101";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000100000";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001010110";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110111";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011110";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001011";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011011";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010011110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000010000001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001001011";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000001111010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001101111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001011001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001011100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001110101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001111100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010000";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001000011";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000000111110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010101010";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010110100";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110001";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000001000011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001110";
    BPixel<="0000000010101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011010100";
    BPixel<="0000000010111010";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001100000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001100000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110000";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111100";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000000";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110010";
    BPixel<="0000000001111100";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000000111111";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000000111011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000000111001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001001111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001001110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000010";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001001011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001110100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001111000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001111011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001110010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001101101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010000010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100111";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000101";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011010";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011011001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011010000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010011";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000010010000";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011000101";
    BPixel<="0000000001111100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001101110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010110110";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000011000011";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011000111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011010000";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011100";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011100000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001000";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011101010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011000001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001000010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010000001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001111000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001110011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001111001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001011000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000111000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001001010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001011";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001100";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001111";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001010010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110100";
    BPixel<="0000000010000111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001111011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001110000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001001101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000110100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010111010";
    BPixel<="0000000010110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110110";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101010";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011100111";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101010";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011011";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001111000";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001000110";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001001001";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001000";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001100";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000101101";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001001101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010111";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001010110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001011100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001011111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010000011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001000111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001111";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011010010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010100";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011011";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011011111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011010011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011010011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000010000111";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001100110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001100100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010100010";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011011110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011010";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011000010";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010111001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010011011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001111010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001111001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001111011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101000";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001100110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000001111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011110";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001011111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001011100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001011101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001011111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001001101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000111000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001000101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000100";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001001110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001010100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000000111111";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000000111010";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001010111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000010000010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000010001000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001111100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001100110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000110010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010101111";
    BPixel<="0000000010100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011100100";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110000";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000010011001";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000010010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001101000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010111101";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010111101";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011000100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001100";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010110";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001100110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000111000";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001001";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001000101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000000111111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001000001";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000101100";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000111000";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001001110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001001001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001110001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000111010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010000010";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001111101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001111000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000001110100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010000000";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010010001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011010111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011010001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011001110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011001001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011100";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010000";
    BPixel<="0000000010001000";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010111110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011011001";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011010001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011001110";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011010000";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011001100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011001101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011000001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010111010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010111000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001111010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010000111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001111010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000101111";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001011011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001110101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001111000";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001000110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001001";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000000111101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001010000";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001101010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001101000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010100001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010101000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000010011101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010110111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010001";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001111001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011001011";
    BPixel<="0000000011000010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001111110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000111110";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011101010";
    BPixel<="0000000010001011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010110001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010110010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010010110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010001100";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010000011";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000010000110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000111101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001110111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001010001";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001001010";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001010110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001000101";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001000000";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000110101";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000110110";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011011";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001110011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010000001";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010000000";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001110001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001010001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000101010";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000010010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000101111";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000110001";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001001";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001111101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001111110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011000001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011000110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010111101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011000111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011010101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000101";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011100000";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110010";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000001001000";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001100111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100010";
    BPixel<="0000000010111101";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000111011";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001101010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011011000";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011011100";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011011111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001011";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011010111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011011100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010011";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010011000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010101111";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000010000100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000001111100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001111000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001000010";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000000111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000101011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000000111000";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101110";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001110010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001001100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000111001";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000000101000";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000101001";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000000111111";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001111101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001000011";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001000000";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001000011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110110";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000111110";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101001";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000010111100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011000000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010100011";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011000010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010101110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010110011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000001001001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011101111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110100";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000001011101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011011";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010100001";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010101001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010101101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010101111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010110000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010100001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010011010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000011";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001111111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001010001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001110";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001000111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001000100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000110000";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000100110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000101010";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000110010";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000000110111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000000111111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001000110";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001001101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000000110010";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000001111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000010110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000000111011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001011010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001110001";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001110101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001111010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001110100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001001111";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010100010";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111110";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000110";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010110";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011100011";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011100011";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011010000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011100100";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011010011";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011010000";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010100101";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000001001011";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000110011";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011001101";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101110";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101101";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011100101";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001101100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000000100101";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000010000001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000010011100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000011000010";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011000100";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000011000010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010110000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010011110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010010100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001101110";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001000000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000000111111";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001111100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010111101";
    GPixel<="0000000001111010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001101110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001110000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001110001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001110011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110110";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001010000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001000111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000000111111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000000110001";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000000111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000010110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000011101";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000011001";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000011001";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000011100";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000100010";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000001";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001110001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001111011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000000111100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001010010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001001001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000011101";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110110";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110101";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110101";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010111001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010110101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000010111011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010011110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010101101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010101101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000010111111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000010101000";
    BPixel<="0000000010011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101011";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001011011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111110";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000100";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111010";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010110100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111000";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101000";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010010011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000001100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000000111111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011110";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001110010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001111010";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001110000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001100011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001000110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001000000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000000111111";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000000111100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000111100";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000000111011";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000000111111";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000000111111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001000000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000000111111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001010011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000001110110";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000001110100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001110000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001111101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001000001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010010000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011001011";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010100110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001110110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000111001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000001000001";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000001000011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010011100";
    BPixel<="0000000010000101";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011011100";
    BPixel<="0000000011001111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110010";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101011";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011110100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110000";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101110";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011010111";
    BPixel<="0000000011001000";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010111010";
    BPixel<="0000000010100011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011011000";
    BPixel<="0000000010110010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000010011011";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000001010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010110";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011000111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010011000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001101111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110011";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001101011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001011111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001011101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001110110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001110011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001101110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001111000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001111010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001111000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001110100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001111010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001111010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001111001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001111000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001110011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001110010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001101111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001111";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001001100";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001001111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001000010";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001000000";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001100000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001111011";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000000110010";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000010000100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000001001100";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001101100";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001111100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010011011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010010110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010011001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010100011";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001100000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000110100";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001001110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010110";
    BPixel<="0000000011000100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011101101";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100101";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110100";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000010001100";
    BPixel<="0000000010000001";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000001100101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000000111010";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001100101";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111111";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000001";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101111";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000111010";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001000100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001010110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001010100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001010110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001100100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001110001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001110000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000001101101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000001101101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000001110101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001110111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111110";
    GPixel<="0000000001001001";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011001001";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011011";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001111110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000010001001";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111000";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110011";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011101101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011101111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111000";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111000";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111001";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110110";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000010000100";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010100011";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011011011";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011010111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010011110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001111101";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001110000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000001110010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001101010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001101001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100010";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011110";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001110";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001001101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010001";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001000110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001001111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010100";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010011100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010101011";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001100010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001111";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011101000";
    BPixel<="0000000010110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011101000";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101000";
    BPixel<="0000000011000010";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001110000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010101111";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010101110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010101111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010111101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001001000";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001100100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001100001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010011";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001001110";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001001101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011110";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001100111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001100111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001100011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000001100100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000001101111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001101010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001011";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111100";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011000110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010011001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010001101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110100";
    GPixel<="0000000010010011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011000101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001101";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010001100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000011001011";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111011";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110001";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110100";
    BPixel<="0000000011010101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000001010000";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011011101";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011010010";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110100";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011010111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010101000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001011101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001101100";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101100";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001101110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001001101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000001110010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000001101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001100101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001100110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001100111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001100111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001100101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001100101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001100111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001011111";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001001111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001011011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111010";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010110010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010110010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010101000";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010101101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010110000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010101100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111110";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001101";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001101100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110011";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011010011";
    BPixel<="0000000011001010";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010101001";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011001011";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010101000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010110101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010101001";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000010111001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000010101001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010100110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000010111100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010110010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010011100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000101";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000001110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000000111001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001110000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001011000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001001100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010011";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001010100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001010111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001010111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001011110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001011101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000001101001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000001101011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001101001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001100110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001100111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001101001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000001110001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001101100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000001110010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001101010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000001110010";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000000111111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000010000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001110100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000100";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010100110";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010111100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011001101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011010110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011010110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011001100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101000";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000000010101";
    GPixel<="0000000000010100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010111110";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110110";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001111001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001011101";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101100";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011010100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011100010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000100";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011010010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011001011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011010101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000100";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010111011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010111001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001010011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000001110110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001101001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001101010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100111";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100101";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100000";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001011111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001011110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001010111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010011";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001010000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001010011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001000111";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000111001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110001";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111011";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010100110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010101000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010100110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000010110101";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000010111001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010100100";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010110110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010110110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010011101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011000010";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000111111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000010010110";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110011";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011110011";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001111111";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000001000001";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010110";
    BPixel<="0000000010001111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010111011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010101110";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000010110001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010100110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010100101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010011011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000000000110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001011100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111000";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010001111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010111";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001010001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011001";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001010000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001010001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001010101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001011010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011000";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001010111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001011111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001011111";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001011110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001011100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001100011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100110";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000001100111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001100110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100111";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001101010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001101110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001110010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001110100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001111000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001011000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001110011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001001";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000010110010";
    GPixel<="0000000010010000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010101001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001011";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010011";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001110";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011011110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011100011";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000010001001";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000001010100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110111";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111100";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111001";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000001011110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001100110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000010100011";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011000101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001011";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011011110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001111";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100100";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011010001";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011000100";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011011001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011001111";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000010001010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001011100";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000110";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011001011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010011111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011001001";
    GPixel<="0000000010100011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001101000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001011001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001100001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001101100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001100100";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001100010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100111";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001100100";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000001100001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100000";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001011110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001011101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001010111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001010101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001010010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001001110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001000111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001100000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001011001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000000110101";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001100";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010100100";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100010";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001111001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110011";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001011111";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001111100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110011";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000000";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010101010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010101111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011000011";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010110110";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010111001";
    BPixel<="0000000010010000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110101";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111001";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000000100011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000010001110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010110001";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000010";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000010";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000011";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010100001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001100000";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000000111100";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000000001110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001100000";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011000011";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010011001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111100";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110001";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011001001";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001011011";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001000110";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001011101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001010001";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001010100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001011110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001011110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011100";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100100";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010100011";
    GPixel<="0000000001101001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000001101010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001100101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001100010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001100110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001101100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001110001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001101011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001010101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000110101";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010010010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101100";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010000";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011011011";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001111000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001100000";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111111";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010111001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111101";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011011011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011010000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010100";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011001110";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011101010";
    BPixel<="0000000010100101";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000001010011";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001110110";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110001";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111001";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101011";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011010000";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011000000";
    GPixel<="0000000010110101";
    BPixel<="0000000001111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110000";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001111";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011010000";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011011011";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000011001110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011010000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011011010";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000011000010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000010000101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000111100";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000001110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001100010";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011011010";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011011000";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011011001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011001011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100100";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000000111110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001100101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000111100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000111100";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001011001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000001100100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001110101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001100111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001011010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000001011101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100011";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001100110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001010111";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001011110";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000010011011";
    GPixel<="0000000001100000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001010101";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010011";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000001010100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001010100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010100";
    GPixel<="0000000001100111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001010111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001000101";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000100110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101010";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000001111001";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010001110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010100110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010101110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010101101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011000101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010110100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001011001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000001000101";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000111100";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000110010";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000110100";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000100011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000111100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000010001101";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011101111";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101100";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110100";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011100010";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011010011";
    BPixel<="0000000011001111";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010101110";
    BPixel<="0000000010100111";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000010011110";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010100101";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010100111";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011011010";
    BPixel<="0000000010111001";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000010011111";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000110101";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010110011";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000010111000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010100011";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010100111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010111110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010100110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000010011101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001001001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001001010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000010111111";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010101000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011001111";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001110010";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001101001";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001000101";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001001111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001010001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000010001111";
    GPixel<="0000000001011100";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010010000";
    GPixel<="0000000001011100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001100000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000001110001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001011111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000001100000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000001101010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001101000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000001101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001100110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000001100010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001010111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000001000001";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000000111101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000001101000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010001001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010110111";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000010001000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010001100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010111011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011010011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010110";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001101";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000100001";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000111000";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001110110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010111000";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000011001101";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000011000111";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011011010";
    BPixel<="0000000010000111";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011101000";
    BPixel<="0000000010100000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000010001111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000001001010";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001110010";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110010";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111010";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111001";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011110011";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001110001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000000111001";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000001010001";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000001000110";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000001010011";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001111110";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010111";
    BPixel<="0000000011000100";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001111000";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000001110010";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011100100";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011000011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010011";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000000";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011111";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011010100";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000001001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111010";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010110011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110111";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001011110";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000001111011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001010100";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001000111";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000000100111";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000000011110";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000000111001";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000000111001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000000111101";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000000";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000001001001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001010000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001000001";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000001001110";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000000110110";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001000110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110010";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000000111111";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000100101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001011101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000000101111";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001010010";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111111";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010001001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010100001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010110110";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010101111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000100111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001100010";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111110";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010110110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010100111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000010111110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000111";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000001010011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000001100001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110000";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110110";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110100";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011101110";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011101010";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110110";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001011001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000001100101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011001100";
    BPixel<="0000000010010000";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110100";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101100";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111001";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001110110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010010011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010101101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010100001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010101101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010101111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111101";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000000110111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001110";
    GPixel<="0000000001101000";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000011";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101100";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101001";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010010010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000010011111";
    GPixel<="0000000001110010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000001011110";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001001011";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001000010";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000100000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001000011";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000000110000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000000110111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000000111111";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000001001011";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000001010000";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000001011010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000000101001";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001000001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010100001";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011000000";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011000000";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000001110001";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010000111";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110000";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110101";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000101";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100001";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010010111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010100110";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011001101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011100000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011011001";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010110";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011100010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011100010";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000010101001";
    GPixel<="0000000010010110";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000110001";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110100";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011100000";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000010110000";
    GPixel<="0000000010101000";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000010011010";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000010011000";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000010011010";
    BPixel<="0000000001111000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011011111";
    BPixel<="0000000011000101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011101110";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110001";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111001";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111011";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111001";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111001";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111001";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110110";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110101";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011110011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000101110";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010110111";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011010111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001111";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011110";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011011";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011011000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001000";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010111111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011011000";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000010100000";
    GPixel<="0000000001111110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001011";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011001001";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011001011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000010100010";
    GPixel<="0000000001111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010001111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010101101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101111";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010100101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000000111111";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001011111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010111000";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000010111000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111000";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010101101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010101010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010101000";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110101";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010000011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000000111010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111000";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111100";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000000";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111011";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000010000110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010011101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101011";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010110101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100100";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000010111111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010111011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111100";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000001001110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010000000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011000110";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011001100";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010101110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010110010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011001010";
    BPixel<="0000000010011000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000101110";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000010001010";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110000";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011110101";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111000";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011110010";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101010";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011100000";
    BPixel<="0000000011010000";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000001010001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000111001";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010110110";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011001010";
    BPixel<="0000000001111101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010100010";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000001010001";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010001010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010100101";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011000000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000110";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000001011010";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000010001100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111010";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010110111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110001";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010101110";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111110";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010100000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000010010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010001101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000010111001";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011000010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010110011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011000101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000001111101";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000000110111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010110101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011000110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011001100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000010000100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110101";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001011";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011001101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011011010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010010";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000001111010";
    GPixel<="0000000001011111";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011000010";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010100";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011011011";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011010001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011011010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011010001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000010010000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010000011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000000110111";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111000";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111001";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110001";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110010";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011100101";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111001";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011100101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000010001000";
    GPixel<="0000000010000100";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001000100";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011001000";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011011011";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011100";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011011110";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011000011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101110";
    BPixel<="0000000010001011";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011010011";
    BPixel<="0000000010000111";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000001001000";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000000010110";
    GPixel<="0000000000000000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000010001110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011001011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011001010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011011000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011011100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011010101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010111011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011010111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010110100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010100011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000101100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111111";
    GPixel<="0000000010011101";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011010011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111010";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111010";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011000111";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010110011";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010101111";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000010110101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010110101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000000101001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011000";
    GPixel<="0000000001111101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011011010";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010101111";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000001";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111001";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000010";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110000";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000001100100";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000010011010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011000010";
    GPixel<="0000000010100000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000010111000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010110110";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101101";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010111101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110000";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011000011";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010011100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000010000001";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001001110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000100100";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000101100";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000000010101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001100100";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011010010";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101011";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101110";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101101";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111001";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011110111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010111";
    BPixel<="0000000011001011";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011000101";
    BPixel<="0000000010111001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011001101";
    BPixel<="0000000011000100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011001111";
    BPixel<="0000000010110111";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000011110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110111";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010101100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111010";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010111001";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000010111110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010110001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000010101001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011011110";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000000101101";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000001111100";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000001110101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001111001";
    GPixel<="0000000001010101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111001";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010100111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000010111010";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010101010";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011000000";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000000110101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111001";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111001";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000010111000";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010111111";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010111001";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000101";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011100100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010110011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110001";
    GPixel<="0000000010010010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010110000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011000010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011001010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010111";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011010100";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011010000";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011100011";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011011011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011101001";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001110011";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000001011111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000001001100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000010001001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000011000110";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011011000";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011010001";
    BPixel<="0000000010000010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011001001";
    BPixel<="0000000010000111";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001100100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001000011";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011101010";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111110";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111000";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110000";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011000001";
    GPixel<="0000000010111101";
    BPixel<="0000000010100000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000001001010";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000100111";
    BPixel<="0000000000000100";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000001001010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000001000100";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000000100100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000000101000";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000010010101";
    GPixel<="0000000010000010";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011100111";
    BPixel<="0000000011010011";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001110011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000001110110";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011100101";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010111";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011010011";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011011100";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010100";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010011";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011010000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010110110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000000";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000010010001";
    GPixel<="0000000001110011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010101010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011011110";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011000011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000010111010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010101110";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010111000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010101011";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010110101";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000000011010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010000101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011010010";
    BPixel<="0000000001111011";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010100100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000010101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011000100";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000010001111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000000100010";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010110001";
    BPixel<="0000000010100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101101";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000000111101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000010";
    GPixel<="0000000001100111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011000010";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010111000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110111";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000010110011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010011010";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000100001";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011011111";
    BPixel<="0000000011010011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110101";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111010";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110100";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111001";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111011";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011110010";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011100011";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000001011011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000001010001";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011001010";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010110100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011001000";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010110110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011011111";
    GPixel<="0000000011001000";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000001011000";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011001100";
    GPixel<="0000000010111110";
    BPixel<="0000000010110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011100110";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000001011111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000110010";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010100001";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010100101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001101";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010110011";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000010011100";
    GPixel<="0000000010001001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000000111011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000110011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010100100";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011001010";
    GPixel<="0000000010101011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000010110111";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000010110111";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000010110110";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000010111101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000010111000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010101010";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011000110";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000010110001";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000000010001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010111001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010101011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011001001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010101110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000110";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011011111";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001111";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011100010";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011011011";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011001111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000000110100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101011";
    GPixel<="0000000010100010";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011100110";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011100110";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000010111000";
    BPixel<="0000000010100001";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010001110";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000010011011";
    BPixel<="0000000010000101";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000010111011";
    BPixel<="0000000010101010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011100111";
    BPixel<="0000000011011001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011110101";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011101011";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111001";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111000";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011101110";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011110101";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110100";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000011000100";
    BPixel<="0000000010110010";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000000101110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110101";
    GPixel<="0000000010110000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011001100";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011001011";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000010111010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011000011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011001011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000010100101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011000100";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000010000001";
    GPixel<="0000000001100110";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000001001000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000000011100";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010010100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011011011";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000010110101";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000010110111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000010011011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101000";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010101111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011010101";
    GPixel<="0000000010110001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011010000";
    GPixel<="0000000010111100";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000010010011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000001011011";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001001100";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000000010111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000001000011";
    BPixel<="0000000000000101";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001001101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000011011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000000111100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011011100";
    BPixel<="0000000011011000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011101011";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011100000";
    BPixel<="0000000010111100";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000001000010";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001000001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101101";
    GPixel<="0000000010100000";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010100001";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000011000101";
    GPixel<="0000000010111001";
    BPixel<="0000000001111111";
    wait for clk_period;
    RPixel<="0000000010001101";
    GPixel<="0000000010000001";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000000110001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000010100100";
    BPixel<="0000000010011000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011101101";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011101110";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111100";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011110111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111110";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111011";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011110111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000010100001";
    GPixel<="0000000010101000";
    BPixel<="0000000010010110";
    wait for clk_period;
    RPixel<="0000000000010100";
    GPixel<="0000000000011000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000000111111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000000011101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000011001";
    GPixel<="0000000000011111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000001100101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000011010010";
    BPixel<="0000000010100111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011111100";
    BPixel<="0000000011010101";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011101111";
    BPixel<="0000000011001110";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000010101111";
    GPixel<="0000000010100010";
    BPixel<="0000000010000000";
    wait for clk_period;
    RPixel<="0000000010001001";
    GPixel<="0000000001111011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000010000110";
    GPixel<="0000000001111100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000010111000";
    BPixel<="0000000010000010";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000001110010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000001011100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001110001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000001001001";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000001100101";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000011010001";
    GPixel<="0000000011001001";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000010101001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011011010";
    GPixel<="0000000010101100";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011000001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000010111011";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000010101000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010101000";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011101010";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000001100110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000001010011";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000010111110";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000010100001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011001010";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010110011";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000010101001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011000101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011001011";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011010000";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011010111";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000000101010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010001100";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011110111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011101010";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011101001";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111010";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111001";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011110111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110001";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011101100";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000001001111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000000100001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111100";
    GPixel<="0000000010011111";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001010";
    BPixel<="0000000001111100";
    wait for clk_period;
    RPixel<="0000000011011110";
    GPixel<="0000000011000010";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011001101";
    BPixel<="0000000010000010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000010111010";
    BPixel<="0000000001110001";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000001110101";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000000100010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000001000110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010101000";
    GPixel<="0000000010111000";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000001011001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000000111111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011010111";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000010111110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000011010010";
    GPixel<="0000000010100001";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000010110100";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000010110011";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000011010110";
    GPixel<="0000000010110001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011001101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000010100100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001101010";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010010001";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001010010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001011101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011111000";
    BPixel<="0000000011000100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011010110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011010110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011101010";
    BPixel<="0000000011001101";
    wait for clk_period;
    RPixel<="0000000010100101";
    GPixel<="0000000011000111";
    BPixel<="0000000010100110";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010001101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010001001";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000001010010";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001100111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001100000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000111101";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000001010110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000000111011";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001100100";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001100110";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000010000011";
    GPixel<="0000000010011100";
    BPixel<="0000000010000110";
    wait for clk_period;
    RPixel<="0000000011000111";
    GPixel<="0000000011011111";
    BPixel<="0000000011001001";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011101100";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011110011";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111001";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110100";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110110";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011110111";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011111010";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111101";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011101100";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001001100";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000000101010";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000000111011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001110111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010000001";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000001110111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010010010";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010000110";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000001111111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010000110";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001101001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001101110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000001010110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000001111001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000010001011";
    GPixel<="0000000010101001";
    BPixel<="0000000010000011";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011110101";
    BPixel<="0000000011001110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011110111";
    BPixel<="0000000011010001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011111111";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001010111";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000001110000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010001001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010010000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000001100011";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000001000101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010111011";
    GPixel<="0000000010110100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011000001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000010101111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010101101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011001011";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011011001";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000001110110";
    GPixel<="0000000001111111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000000110110";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000001101010";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000001101100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010000101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000001011001";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000000110010";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000001000000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000001010001";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000001101000";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000001010010";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000000101001";
    BPixel<="0000000000000110";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000001101111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110011";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110110";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110000";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011110011";
    GPixel<="0000000011110011";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011110011";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111001";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111010";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111010";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011101001";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111010";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111000";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011001101";
    GPixel<="0000000011011101";
    BPixel<="0000000010110110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001011010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000000101011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001000110";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000001101110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000010101001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010100110";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010100001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001111011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010100010";
    BPixel<="0000000001111101";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001011110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000010100";
    GPixel<="0000000000111000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000010000111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000010110101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000010111111";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000010110011";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000010110011";
    GPixel<="0000000010011001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000001010111";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000001110";
    GPixel<="0000000000101000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000010110100";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010101010";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001110101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001101110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000001110";
    GPixel<="0000000001000110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000010101010";
    GPixel<="0000000011010101";
    BPixel<="0000000011000001";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011001111";
    GPixel<="0000000011101111";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000001101001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001011110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010001111";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010000101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010010001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010001011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010010011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010001100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001110010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010000001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010010000";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000001110111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000001000";
    GPixel<="0000000001001101";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000001101110";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000001111001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000000101";
    GPixel<="0000000000110111";
    BPixel<="0000000000000010";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010110010";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011101100";
    BPixel<="0000000011010111";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000011011101";
    BPixel<="0000000011011010";
    wait for clk_period;
    RPixel<="0000000010111010";
    GPixel<="0000000011000110";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000010111001";
    GPixel<="0000000011001010";
    BPixel<="0000000011000000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000011010101";
    BPixel<="0000000011000111";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011100101";
    BPixel<="0000000011011000";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011110100";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011111101";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011000110";
    GPixel<="0000000011011100";
    BPixel<="0000000011000101";
    wait for clk_period;
    RPixel<="0000000010001100";
    GPixel<="0000000010101001";
    BPixel<="0000000010001101";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000001110101";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000001010101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000001001100";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000001010100";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000001011100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001001110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001011000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000001011101";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001011111";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000011000";
    GPixel<="0000000001011011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000001011011";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000000011011";
    GPixel<="0000000001101000";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000001101110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000000010001";
    GPixel<="0000000001100000";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010000001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010001011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010001000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010001001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010001001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010010000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010001111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010010110";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010000111";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010010000";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010000110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000001100000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011010100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000010010111";
    GPixel<="0000000011001101";
    BPixel<="0000000010110011";
    wait for clk_period;
    RPixel<="0000000000000010";
    GPixel<="0000000001000001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000001111110";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010010100";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010001100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010100010";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000001111110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000001000100";
    BPixel<="0000000000000001";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000000101111";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000001001001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000001010000";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000011000";
    GPixel<="0000000000101101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000001000";
    GPixel<="0000000000110001";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000001110100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010010011";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010000101";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010000111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010001010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010001100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010100001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001111100";
    GPixel<="0000000010111010";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010010101";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001011001";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000001001111";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000010010011";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111011";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111101";
    BPixel<="0000000011110000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110100";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111100";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111100";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000010011010";
    GPixel<="0000000010101000";
    BPixel<="0000000010011001";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000000101100";
    BPixel<="0000000000001111";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001100001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000001011010";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000000000100";
    GPixel<="0000000001000000";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010101001";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010011111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010010000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000010001010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010001010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010001010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000001111111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000001101011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000001011011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000001011101";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000001100100";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001101010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000010110";
    GPixel<="0000000001010100";
    BPixel<="0000000000010001";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010011000";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010101011";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010001001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010000001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000010100";
    GPixel<="0000000001010111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010000011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010011000";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001101011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010101101";
    BPixel<="0000000001110010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000001111110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010000100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010010011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010001000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010001101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010010100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010000110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010000111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010001000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000010101";
    GPixel<="0000000001100101";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000011000010";
    BPixel<="0000000001111001";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001110000";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000000110";
    GPixel<="0000000001011001";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010001000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010011011";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010010000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010010010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010011110";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010010111";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010100100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010100111";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010010001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001101111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000000010110";
    GPixel<="0000000001011101";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001100110";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000001110100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000011010010";
    BPixel<="0000000010111000";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011111011";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011110100";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111100";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111001";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011101101";
    BPixel<="0000000011100101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011101011";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000010010010";
    GPixel<="0000000010111000";
    BPixel<="0000000010011111";
    wait for clk_period;
    RPixel<="0000000000010001";
    GPixel<="0000000001001000";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000001111011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010010001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010100111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010101101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010100110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010011110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010011110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010011011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110000";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101111";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010100001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010100010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010100000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010000111";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000011000";
    GPixel<="0000000001101010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000001110";
    GPixel<="0000000001100000";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001110000";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010001110";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010010000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010000001";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010010100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010011110";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000011011";
    GPixel<="0000000001111101";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010001100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010000111";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010010100";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010011001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000001001011";
    BPixel<="0000000000000011";
    wait for clk_period;
    RPixel<="0000000000010111";
    GPixel<="0000000001100100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000001010101";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000001100110";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000001111100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010011010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010101110";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000001110111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000000111";
    GPixel<="0000000001010100";
    BPixel<="0000000000001110";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001110101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010010101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010001111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010000101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010001011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010010001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010010110";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010010111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010010100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010010100";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000010000111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010111001";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010010101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010001001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000001011011";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000001101011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000001010000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000001001111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111100";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111011";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000001010111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001011010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000000101001";
    BPixel<="0000000000001010";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000010100100";
    BPixel<="0000000001110011";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010011101";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010100001";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010011001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000010001100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000010010000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010010010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010001111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010001010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010000101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010000111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010001010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010000100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010011100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010001010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010000000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000001101100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010011111";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010100110";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010000011";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000001111101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000001001110";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000011001";
    GPixel<="0000000001101100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000001101";
    GPixel<="0000000001100100";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000010000101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010010001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010000100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010010110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010001000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010001101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000010000001";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010010010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010001100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000001100001";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000001111110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010011100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010101101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010100110";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010100110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010100001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010101101";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010100011";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010010110";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000001111101";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000010010";
    GPixel<="0000000001000001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010000111";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111010";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011101101";
    BPixel<="0000000011100100";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111001";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000010100011";
    BPixel<="0000000010001001";
    wait for clk_period;
    RPixel<="0000000000010101";
    GPixel<="0000000001000001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010000010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000010110100";
    BPixel<="0000000001110111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010101010";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010100010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010011000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010011001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101110";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010011011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010100010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010101001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010000101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010010101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010100001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010100110";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010011100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000001010010";
    BPixel<="0000000000001001";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001110101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010100000";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010000100";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010001100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010011001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010001100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010000111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010001011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010100000";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010001011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000001100110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010001101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010001110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010101001";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010001001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001111100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010100010";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010001101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010000111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000001110111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010001101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010001001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010000111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010001010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010011011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010110100";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000010101110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010000000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000010010110";
    GPixel<="0000000010111111";
    BPixel<="0000000010010011";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000001011111";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000001000111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001110010";
    GPixel<="0000000001111000";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011011111";
    BPixel<="0000000011011110";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000001001010";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000001010101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000010010010";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000001100101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010101110";
    BPixel<="0000000001100110";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000011000000";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010011011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010000";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010010000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000010001110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000010001110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010001111";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010010010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010010011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010011100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010000110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000010000010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010001000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001111101";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001111110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010101110";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010010101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010001011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000010110";
    GPixel<="0000000001101101";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000011011";
    GPixel<="0000000001110101";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010101010";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010011000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010001010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010011100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000010000110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010010101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010000110";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010010010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001111000";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000010001";
    GPixel<="0000000001101001";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010010000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010011101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010010000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001111011";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010010001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010100";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010100011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010100000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010011111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010011110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010101011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010100110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010010111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000010111011";
    BPixel<="0000000001111010";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000001111001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000011000";
    GPixel<="0000000001000010";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000011001110";
    GPixel<="0000000011101000";
    BPixel<="0000000011001101";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111110";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111001";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011111111";
    BPixel<="0000000011100111";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000001110000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010000100";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010100110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010010000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010011110";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010100111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010101111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010101010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010101011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010100100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010011101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010011001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010011010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010100110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010100000";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000001111010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001111001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010110101";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010010000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000001001";
    GPixel<="0000000001100011";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000001111110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001111111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010011010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000010000011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100011";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000010000101";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010010110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000001100111";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001111010";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010001000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010100101";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010100110";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000000011011";
    GPixel<="0000000001110101";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000011001";
    GPixel<="0000000001110101";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000001111000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010010011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010011100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010001";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010010010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010010000";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010001100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010001100";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010010011";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010011000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000011000001";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010011011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001101011";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001111111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000010111110";
    GPixel<="0000000011100010";
    BPixel<="0000000010111100";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000011010000";
    BPixel<="0000000010111010";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000010111110";
    BPixel<="0000000010110100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111010";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111010";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111011";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010000101";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000001001111";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000001010000";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010101110";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010110001";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010110011";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010101010";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010011110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010100";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010010100";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010010100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010010011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010000101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010100100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010000001";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000010111";
    GPixel<="0000000001110010";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001111110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010101110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010001101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010001100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001111000";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000001111110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010001001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010000010";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010011010";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010001110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000001111000";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010011111";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000001100100";
    BPixel<="0000000000011010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010010011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010100010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000001110";
    GPixel<="0000000001101001";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010011001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010011011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010101000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010011010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110010";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101110";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010100111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010100110";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100111";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010101001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010100010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010100011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010100111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010100011";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010101010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010101000";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000000111010";
    BPixel<="0000000000001011";
    wait for clk_period;
    RPixel<="0000000011001011";
    GPixel<="0000000011100110";
    BPixel<="0000000011000111";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011101110";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111010";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010000110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001100110";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000010111000";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010100011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010101100";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010110010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010101111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010110000";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010101111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010101100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010100001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000010011111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010100110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000010011101";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100100";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010011100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010100100";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110011";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010100111";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101000";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000001111111";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000001111110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010000010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000001101011";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010011101";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010001100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010001111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010001110";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010000101";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000001011";
    GPixel<="0000000001100010";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000001111001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010001010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010010001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010100010";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000001010011";
    BPixel<="0000000000000111";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000001110101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010010110";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010100101";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010010111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010010100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010010000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010001101";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000010001001";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000010000111";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000100011";
    GPixel<="0000000010001011";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010010111";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010100101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010101110";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010101110";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010101011";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001110100";
    GPixel<="0000000010110110";
    BPixel<="0000000001101111";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000001101100";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000011010101";
    BPixel<="0000000010101011";
    wait for clk_period;
    RPixel<="0000000011100110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011111000";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011101001";
    BPixel<="0000000011011111";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111101";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111111";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011110111";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111000";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011110101";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011100101";
    GPixel<="0000000011110011";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011011001";
    GPixel<="0000000011111001";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000011011000";
    GPixel<="0000000011111101";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000010100100";
    GPixel<="0000000011010100";
    BPixel<="0000000010100010";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000001111000";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000001100100";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010000101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010000100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000010000000";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000010000010";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000010000100";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000010001000";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000100001";
    GPixel<="0000000010001010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000010000111";
    BPixel<="0000000000100101";
    wait for clk_period;
    RPixel<="0000000000010100";
    GPixel<="0000000001111100";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000001110";
    GPixel<="0000000001110011";
    BPixel<="0000000000010011";
    wait for clk_period;
    RPixel<="0000000000001011";
    GPixel<="0000000001101011";
    BPixel<="0000000000010010";
    wait for clk_period;
    RPixel<="0000000000010110";
    GPixel<="0000000001110101";
    BPixel<="0000000000100001";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010000011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000010000000";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010100010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010100111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000011001";
    GPixel<="0000000001101101";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000001100011";
    BPixel<="0000000000011000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010101011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010010011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000100100";
    GPixel<="0000000001110110";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001111011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000001011111";
    BPixel<="0000000000011001";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010000000";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010011000";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010001111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001111110";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000000010001";
    GPixel<="0000000001101001";
    BPixel<="0000000000011101";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001110110";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010011000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010100011";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010100110";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010101000";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010100111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010101010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010101100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010101010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010100001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010100111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010101010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010101011";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000010101010";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010101011";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010111010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010101011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010010100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000001010010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011110100";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111101";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000010111000";
    GPixel<="0000000011010000";
    BPixel<="0000000010111000";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000001010111";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000010101110";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010110101";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010100101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010101101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010111011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010110000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100100";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010101010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010101011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010100101";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010100001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010011101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010001101";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000001110100";
    BPixel<="0000000000100110";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000001100111";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010001001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010100001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000000011101";
    GPixel<="0000000001101101";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000001101";
    GPixel<="0000000001011101";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001111001";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000001111100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010011111";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010011101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000001110010";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010001111";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010000010";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000001110010";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000001111110";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000010000010";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010001110";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010100111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110001";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110100";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010111001";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010111011";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010111001";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010110110";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010110010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010011111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010101100";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010001100";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000001101011";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000001101110";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001110111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010010010";
    BPixel<="0000000001101110";
    wait for clk_period;
    RPixel<="0000000010100110";
    GPixel<="0000000011001001";
    BPixel<="0000000010101011";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111101";
    BPixel<="0000000011101011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111000";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011111010";
    GPixel<="0000000011111000";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011111001";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011100100";
    GPixel<="0000000011111111";
    BPixel<="0000000011100000";
    wait for clk_period;
    RPixel<="0000000010011101";
    GPixel<="0000000010111101";
    BPixel<="0000000010010110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000001110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000001100110";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000001110111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010011010";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000010110000";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010101100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010110001";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010101100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010101010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010101110";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010101001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010011111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010001110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010000000";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010001111";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000001100010";
    BPixel<="0000000000010000";
    wait for clk_period;
    RPixel<="0000000000010011";
    GPixel<="0000000001100100";
    BPixel<="0000000000010101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010011000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010010101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010010011";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000001110011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000010101";
    GPixel<="0000000001100000";
    BPixel<="0000000000011011";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010011110";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000001111101";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000000001";
    GPixel<="0000000001010101";
    BPixel<="0000000000001000";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010000111";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010100101";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010100010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010011111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010100101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101011";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010100111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010100111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100111";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010101011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010110000";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010110100";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010110011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010101111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000011000001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010101111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010110000";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010101111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000010101111";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000001011000";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000010010011";
    GPixel<="0000000010101101";
    BPixel<="0000000010010010";
    wait for clk_period;
    RPixel<="0000000011110110";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000001111101";
    GPixel<="0000000010011010";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000001100010";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010100110";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010100110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000011000101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010111101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010111011";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010111001";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110111";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101000";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010100110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010100110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101011";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010101000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010100010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010100011";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010100011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010101101";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010011000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000001011";
    GPixel<="0000000001100010";
    BPixel<="0000000000010100";
    wait for clk_period;
    RPixel<="0000000000011010";
    GPixel<="0000000001100111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010001001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001101001";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010000111";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010010010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010001111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001111001";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000000000000";
    GPixel<="0000000001001101";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010001010";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010001101";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010011010";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010110000";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010110100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000011001101";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010110101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010101111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010101101";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010111111";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010110010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010101000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010101010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010101101";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010101010";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000010100000";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010000100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000001011100";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001110000";
    GPixel<="0000000010011010";
    BPixel<="0000000001101100";
    wait for clk_period;
    RPixel<="0000000011100010";
    GPixel<="0000000011111111";
    BPixel<="0000000011011101";
    wait for clk_period;
    RPixel<="0000000011101111";
    GPixel<="0000000011111111";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011111001";
    BPixel<="0000000011100011";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011110000";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011011011";
    GPixel<="0000000011101000";
    BPixel<="0000000011010110";
    wait for clk_period;
    RPixel<="0000000011101011";
    GPixel<="0000000011111111";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011100001";
    GPixel<="0000000011111111";
    BPixel<="0000000011011100";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000001110001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000001110001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010011100";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001111000";
    GPixel<="0000000010111011";
    BPixel<="0000000001110100";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010100101";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010101001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010101101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010111100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010111000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010101011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101010";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010110111";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010110110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010110111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010110111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010110110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010101110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010011111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010100010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010011011";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010000110";
    BPixel<="0000000000100011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010010100";
    BPixel<="0000000000110011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010010111";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000001111101";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010001101";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000101001";
    GPixel<="0000000010000001";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000011000";
    GPixel<="0000000001110000";
    BPixel<="0000000000011100";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001111011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001110001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000001111110";
    BPixel<="0000000000110010";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001110010";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000001101010";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000001000";
    GPixel<="0000000001011001";
    BPixel<="0000000000001101";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010000101";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001000010";
    GPixel<="0000000010100001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010100110";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101010";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010100001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010101001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010101011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101011";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010101000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010100111";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111101";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010111010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010110000";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010100011";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010100001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010101011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010101110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000011000001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010101010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000010110100";
    BPixel<="0000000001101000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000001110001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000010001001";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001111100";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000001110000";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000010111100";
    BPixel<="0000000001110000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010101110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010110011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010101110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000011000011";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010110001";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010110010";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010110010";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010110001";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010101110";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101110";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010110100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010110110";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010101101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010101010";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010101001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010101100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010101100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010101010";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110000";
    GPixel<="0000000010101100";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010100101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010101011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010100010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010011110";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010100011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010100010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000000010001";
    GPixel<="0000000001100100";
    BPixel<="0000000000010110";
    wait for clk_period;
    RPixel<="0000000000001010";
    GPixel<="0000000001011000";
    BPixel<="0000000000001100";
    wait for clk_period;
    RPixel<="0000000000100000";
    GPixel<="0000000001110001";
    BPixel<="0000000000100100";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000001111011";
    BPixel<="0000000000101011";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010000001";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010011001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010010001";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010101101";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010100001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010101110";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010111111";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010101111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010010111";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100011";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010101001";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010110000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010110101";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010111000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000011001011";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010111101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010111001";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010111101";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010111100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010101110";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010101100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010101101";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000010101100";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000001110001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000001110011";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011101101";
    GPixel<="0000000011111111";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011110011";
    wait for clk_period;
    RPixel<="0000000011010111";
    GPixel<="0000000011101011";
    BPixel<="0000000011010000";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000011001110";
    BPixel<="0000000010100111";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000001101000";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000001110001";
    GPixel<="0000000010101101";
    BPixel<="0000000001101101";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010101101";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010110110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010111110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010111111";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010111011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000011000001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000011001001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000011001001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000011000001";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010110110";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000011001000";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000011000101";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000011000000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010111100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010111010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111000";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010110110";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000011000100";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101111";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111010";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010111101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111100";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000011000101";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010111010";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010101111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010110110";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010111000";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010101001";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010010010";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010000110";
    BPixel<="0000000000110101";
    wait for clk_period;
    RPixel<="0000000000011100";
    GPixel<="0000000001101111";
    BPixel<="0000000000011111";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000001111001";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010101010";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100001";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010100000";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010100101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000010100101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101010";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000010101100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010101000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000010101001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010101100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000101111";
    GPixel<="0000000010101100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010101011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010110001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010111101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010111110";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010111011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000010111011";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000010111001";
    BPixel<="0000000001101010";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000010110010";
    BPixel<="0000000001101001";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010101001";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010100010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010111100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010110101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010110110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010110001";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000010110000";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000001100101";
    BPixel<="0000000000110000";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000001111111";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010000111";
    BPixel<="0000000001100111";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000001100010";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010100001";
    BPixel<="0000000001011100";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000010110100";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000011000000";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010100100";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000001111010";
    BPixel<="0000000000101001";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000001111101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000001100100";
    BPixel<="0000000000101010";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001011000";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000001110000";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010100000";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000010111110";
    BPixel<="0000000001100011";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100111";
    BPixel<="0000000000111000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010101111";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010101100";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010101001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010101010";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000010101011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000101101";
    GPixel<="0000000010101011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000000101100";
    GPixel<="0000000010101001";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000101000";
    GPixel<="0000000010100010";
    BPixel<="0000000000111101";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010110010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000010101010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000110001";
    GPixel<="0000000010100000";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010101000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000000111000";
    GPixel<="0000000010011111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010100101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000010000011";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010011001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010101110";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101001";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101100";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010100100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000011000101";
    BPixel<="0000000001100010";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111000";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110010";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101101";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000011000000";
    BPixel<="0000000001010100";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010101110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000011001010";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010110000";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010110000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010101101";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010101110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010110101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010111100";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010111110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000010111111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000011000010";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000011000100";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111110";
    BPixel<="0000000000111011";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111100";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000011000011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000011000001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010111101";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010111110";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010110111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010110011";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010001011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000001101111";
    BPixel<="0000000000110100";
    wait for clk_period;
    RPixel<="0000000000110011";
    GPixel<="0000000001010110";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111100";
    GPixel<="0000000011111110";
    BPixel<="0000000011111001";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111101";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111101";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011111000";
    GPixel<="0000000011111111";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000010110110";
    GPixel<="0000000011001101";
    BPixel<="0000000010110001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000001101010";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000000100110";
    GPixel<="0000000001011001";
    BPixel<="0000000000010111";
    wait for clk_period;
    RPixel<="0000000000001100";
    GPixel<="0000000001001011";
    BPixel<="0000000000000000";
    wait for clk_period;
    RPixel<="0000000001111011";
    GPixel<="0000000011000111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010110001";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010110111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010111100";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001100010";
    GPixel<="0000000010111011";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010111011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010111011";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010111100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000010111110";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010111111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011110";
    GPixel<="0000000011000010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010011";
    GPixel<="0000000010111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010110111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010110111";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010110100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010110011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010111001";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010011100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010011011";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000011110";
    GPixel<="0000000010000110";
    BPixel<="0000000000110001";
    wait for clk_period;
    RPixel<="0000000000011111";
    GPixel<="0000000010001001";
    BPixel<="0000000000101111";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010110100";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110001";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010100111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010101100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000000111101";
    GPixel<="0000000010101001";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010110001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010110011";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000000111100";
    GPixel<="0000000010110001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010111011";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000000111011";
    GPixel<="0000000010101111";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110101";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001010111";
    GPixel<="0000000010111101";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010110100";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001011000";
    GPixel<="0000000010110010";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010101001";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000010101111";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000010000100";
    GPixel<="0000000011000001";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001110110";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000000100101";
    GPixel<="0000000001000111";
    BPixel<="0000000000100010";
    wait for clk_period;
    RPixel<="0000000001110111";
    GPixel<="0000000010001101";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000011001000";
    GPixel<="0000000011011001";
    BPixel<="0000000011000110";
    wait for clk_period;
    RPixel<="0000000011101001";
    GPixel<="0000000011111100";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000011011101";
    GPixel<="0000000011111000";
    BPixel<="0000000011011001";
    wait for clk_period;
    RPixel<="0000000010011110";
    GPixel<="0000000011000101";
    BPixel<="0000000010011000";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000001110110";
    BPixel<="0000000000111111";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010010011";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000010101100";
    BPixel<="0000000001101011";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000010011100";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000000110100";
    GPixel<="0000000001011001";
    BPixel<="0000000000101101";
    wait for clk_period;
    RPixel<="0000000010001010";
    GPixel<="0000000010100101";
    BPixel<="0000000010000100";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011101100";
    GPixel<="0000000011111011";
    BPixel<="0000000011100110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000011000111";
    BPixel<="0000000010100111";
    wait for clk_period;
    RPixel<="0000000000100111";
    GPixel<="0000000001000111";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000010000111";
    GPixel<="0000000010101101";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000001111111";
    GPixel<="0000000010101010";
    BPixel<="0000000001110101";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000001101001";
    BPixel<="0000000000110111";
    wait for clk_period;
    RPixel<="0000000010011001";
    GPixel<="0000000010110111";
    BPixel<="0000000010010001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011111101";
    BPixel<="0000000011110010";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011110111";
    BPixel<="0000000011110101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011000100";
    GPixel<="0000000011010010";
    BPixel<="0000000011000001";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000001101001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000101011";
    GPixel<="0000000001010101";
    BPixel<="0000000000100111";
    wait for clk_period;
    RPixel<="0000000010000101";
    GPixel<="0000000010111101";
    BPixel<="0000000001111110";
    wait for clk_period;
    RPixel<="0000000001101111";
    GPixel<="0000000010110111";
    BPixel<="0000000001100101";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010110101";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010101000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010111010";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000011000100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001000001";
    GPixel<="0000000010110011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010111101";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110101";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110111";
    BPixel<="0000000001010010";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010110110";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000000010111";
    GPixel<="0000000010000110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000000100010";
    GPixel<="0000000010001110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000000110111";
    GPixel<="0000000010100011";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000000110101";
    GPixel<="0000000010100010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010111100";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010110110";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010111001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010111001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010111000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010111001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001011100";
    GPixel<="0000000010111110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011111";
    GPixel<="0000000010111100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010111100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010111011";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010111010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000010111010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000010111011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010111001";
    BPixel<="0000000000111110";
    wait for clk_period;
    RPixel<="0000000001110011";
    GPixel<="0000000011001000";
    BPixel<="0000000001010011";
    wait for clk_period;
    RPixel<="0000000001100110";
    GPixel<="0000000010110011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010100111";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000001111001";
    BPixel<="0000000000110110";
    wait for clk_period;
    RPixel<="0000000010101110";
    GPixel<="0000000011010010";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000011100000";
    GPixel<="0000000011110111";
    BPixel<="0000000011011011";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011100011";
    GPixel<="0000000011111010";
    BPixel<="0000000011011110";
    wait for clk_period;
    RPixel<="0000000010000000";
    GPixel<="0000000010100100";
    BPixel<="0000000001110110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010000011";
    BPixel<="0000000001000000";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000010110101";
    BPixel<="0000000001011110";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010110010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010110110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010110101";
    BPixel<="0000000000111010";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010111010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010111011";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010111100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010111101";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010111011";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010111100";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001011101";
    GPixel<="0000000010111010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010111011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010101";
    GPixel<="0000000010111000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010010";
    GPixel<="0000000010111001";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010111000";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111001";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010111001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010111010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110110";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010111110";
    BPixel<="0000000001011011";
    wait for clk_period;
    RPixel<="0000000000111001";
    GPixel<="0000000010100110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000000111110";
    GPixel<="0000000010101010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000010010110";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000000001111";
    GPixel<="0000000001111110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010101110";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110100";
    BPixel<="0000000001010001";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110010";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010111010";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110111";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111010";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111011";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110101";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000011000100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010111100";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001001101";
    GPixel<="0000000010111000";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000010110000";
    BPixel<="0000000001001011";
    wait for clk_period;
    RPixel<="0000000001010000";
    GPixel<="0000000010101010";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001100100";
    GPixel<="0000000010111000";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001101011";
    GPixel<="0000000010110011";
    BPixel<="0000000001100001";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000001101100";
    BPixel<="0000000000101110";
    wait for clk_period;
    RPixel<="0000000001001110";
    GPixel<="0000000001110101";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000011000011";
    GPixel<="0000000011011101";
    BPixel<="0000000011000000";
    wait for clk_period;
    RPixel<="0000000011110111";
    GPixel<="0000000011111111";
    BPixel<="0000000011110110";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011110000";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111100";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111100";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101111";
    wait for clk_period;
    RPixel<="0000000011100111";
    GPixel<="0000000011111111";
    BPixel<="0000000011100001";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000010001111";
    BPixel<="0000000001100000";
    wait for clk_period;
    RPixel<="0000000001101110";
    GPixel<="0000000010010110";
    BPixel<="0000000001100100";
    wait for clk_period;
    RPixel<="0000000001101001";
    GPixel<="0000000010001101";
    BPixel<="0000000001011111";
    wait for clk_period;
    RPixel<="0000000000110110";
    GPixel<="0000000001010101";
    BPixel<="0000000000101100";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011111111";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011101000";
    GPixel<="0000000011110111";
    BPixel<="0000000011100010";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011110111";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111110";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111101";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111110";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110000";
    GPixel<="0000000011111101";
    BPixel<="0000000011101001";
    wait for clk_period;
    RPixel<="0000000011110100";
    GPixel<="0000000011111111";
    BPixel<="0000000011101100";
    wait for clk_period;
    RPixel<="0000000001011010";
    GPixel<="0000000001111001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000001101000";
    BPixel<="0000000000111100";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010000001";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000010101100";
    GPixel<="0000000011010000";
    BPixel<="0000000010100100";
    wait for clk_period;
    RPixel<="0000000011101110";
    GPixel<="0000000011111111";
    BPixel<="0000000011101000";
    wait for clk_period;
    RPixel<="0000000011011100";
    GPixel<="0000000011101110";
    BPixel<="0000000011011000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011110101";
    GPixel<="0000000011110011";
    BPixel<="0000000011110100";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011101010";
    GPixel<="0000000011101010";
    BPixel<="0000000011101010";
    wait for clk_period;
    RPixel<="0000000011110010";
    GPixel<="0000000011111111";
    BPixel<="0000000011110001";
    wait for clk_period;
    RPixel<="0000000011110001";
    GPixel<="0000000011111111";
    BPixel<="0000000011101101";
    wait for clk_period;
    RPixel<="0000000010110111";
    GPixel<="0000000011011110";
    BPixel<="0000000010110010";
    wait for clk_period;
    RPixel<="0000000000110010";
    GPixel<="0000000001100110";
    BPixel<="0000000000101000";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010010100";
    BPixel<="0000000001000010";
    wait for clk_period;
    RPixel<="0000000001100011";
    GPixel<="0000000010110111";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001100001";
    GPixel<="0000000010111011";
    BPixel<="0000000001011001";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010111011";
    BPixel<="0000000001010110";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110111";
    BPixel<="0000000001001101";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010110000";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010111001";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001000100";
    GPixel<="0000000010110110";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001000011";
    GPixel<="0000000010110011";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110011";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001100";
    GPixel<="0000000010110101";
    BPixel<="0000000001010000";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010101111";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001000110";
    GPixel<="0000000010110010";
    BPixel<="0000000001001111";
    wait for clk_period;
    RPixel<="0000000000111111";
    GPixel<="0000000010101101";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000000001101";
    GPixel<="0000000001111100";
    BPixel<="0000000000011110";
    wait for clk_period;
    RPixel<="0000000000101110";
    GPixel<="0000000010011010";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001000000";
    GPixel<="0000000010101100";
    BPixel<="0000000001010111";
    wait for clk_period;
    RPixel<="0000000000111010";
    GPixel<="0000000010100111";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010111101";
    BPixel<="0000000001011010";
    wait for clk_period;
    RPixel<="0000000001000101";
    GPixel<="0000000010110101";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001000111";
    GPixel<="0000000010111000";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010110111";
    BPixel<="0000000001001110";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001100";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111000";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001000";
    GPixel<="0000000010111001";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001010";
    GPixel<="0000000010111010";
    BPixel<="0000000001001010";
    wait for clk_period;
    RPixel<="0000000001001001";
    GPixel<="0000000010111001";
    BPixel<="0000000001001001";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111001";
    BPixel<="0000000001001000";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010110111";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001001011";
    GPixel<="0000000010111000";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001001111";
    GPixel<="0000000010110111";
    BPixel<="0000000001000110";
    wait for clk_period;
    RPixel<="0000000001010001";
    GPixel<="0000000010111000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001010100";
    GPixel<="0000000010110111";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001010110";
    GPixel<="0000000010111000";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001011011";
    GPixel<="0000000010111000";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100000";
    GPixel<="0000000010111011";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010111100";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001100111";
    GPixel<="0000000010111111";
    BPixel<="0000000001000101";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010111101";
    BPixel<="0000000001000100";
    wait for clk_period;
    RPixel<="0000000001101000";
    GPixel<="0000000010111100";
    BPixel<="0000000001000011";
    wait for clk_period;
    RPixel<="0000000001100101";
    GPixel<="0000000010111010";
    BPixel<="0000000001000001";
    wait for clk_period;
    RPixel<="0000000001101010";
    GPixel<="0000000011000010";
    BPixel<="0000000001000111";
    wait for clk_period;
    RPixel<="0000000001011001";
    GPixel<="0000000010101110";
    BPixel<="0000000000111001";
    wait for clk_period;
    RPixel<="0000000001110101";
    GPixel<="0000000011000010";
    BPixel<="0000000001011000";
    wait for clk_period;
    RPixel<="0000000001101100";
    GPixel<="0000000010101100";
    BPixel<="0000000001010101";
    wait for clk_period;
    RPixel<="0000000001101101";
    GPixel<="0000000010100000";
    BPixel<="0000000001011101";
    wait for clk_period;
    RPixel<="0000000000101010";
    GPixel<="0000000001001110";
    BPixel<="0000000000100000";
    wait for clk_period;
    RPixel<="0000000011010011";
    GPixel<="0000000011101010";
    BPixel<="0000000011001110";
    wait for clk_period;
    RPixel<="0000000011111001";
    GPixel<="0000000011111111";
    BPixel<="0000000011111000";
    wait for clk_period;
    RPixel<="0000000011111011";
    GPixel<="0000000011111100";
    BPixel<="0000000011111110";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111011";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111100";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111110";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111110";
    GPixel<="0000000011111111";
    BPixel<="0000000011111011";
    wait for clk_period;
    RPixel<="0000000011111101";
    GPixel<="0000000011111111";
    BPixel<="0000000011111010";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111101";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;
    RPixel<="0000000011111111";
    GPixel<="0000000011111111";
    BPixel<="0000000011111111";
    wait for clk_period;



      -- insert stimulus here 

      wait;
   end process;

END;
